`timescale 100ps / 100ps
//
`default_nettype none

module Top (
    input wire sys_clk,  // 27 MHz
    input wire sys_rst_n,
    output reg [5:0] led,
    input wire uart_rx,
    output wire uart_tx,
    input wire btn1,

    // magic ports for PSRAM to be inferred
    output wire [ 1:0] O_psram_ck,
    output wire [ 1:0] O_psram_ck_n,
    inout  wire [ 1:0] IO_psram_rwds,
    inout  wire [15:0] IO_psram_dq,
    output wire [ 1:0] O_psram_reset_n,
    output wire [ 1:0] O_psram_cs_n,

    // flash
    output reg  flash_clk,
    input  wire flash_miso,
    output reg  flash_mosi,
    output reg  flash_cs
);

  // ----------------------------------------------------------
  // -- Gowin_rPLLs
  // ----------------------------------------------------------
  wire rpll_clkin = sys_clk;
  wire rpll_lock;
  wire rpll_clkout;
  wire rpll_clkoutp;
  wire rpll_clkoutd;

  Gowin_rPLL rpll (
      .clkin(rpll_clkin),  // 27 MHz
      .lock(rpll_lock),
      .clkout(rpll_clkout),  // 81 MHz
      .clkoutp(rpll_clkoutp),  // clkout 81 MHz 90 degrees phased
      .clkoutd(rpll_clkoutd)  // clkout / 4 = 20.25 MHz (IPUG943-1.2E page 15)
  );

  // ----------------------------------------------------------
  // -- PSRAM_Memory_Interface_HS_V2_Top
  // ----------------------------------------------------------
  wire br_clk_d = rpll_clkoutd;
  wire br_pll_lock = rpll_lock;
  wire br_memory_clk = rpll_clkout;
  wire br_memory_clk_p = rpll_clkoutp;
  wire br_clk_out;
  wire rst_n = sys_rst_n;
  wire [63:0] br_wr_data;
  wire [63:0] br_rd_data;
  wire br_rd_data_valid;
  wire [20:0] br_addr;
  wire br_cmd;
  wire br_cmd_en;
  wire br_init_calib;
  wire [7:0] br_data_mask;

  PSRAM_Memory_Interface_HS_V2_Top br (
      .rst_n(rst_n),
      .clk_d(br_clk_d),
      .memory_clk(br_memory_clk),
      .memory_clk_p(br_memory_clk_p),
      .clk_out(br_clk_out),  // memory_clk / 2
      .pll_lock(br_pll_lock),
      .init_calib(br_init_calib),

      .cmd(br_cmd),
      .cmd_en(br_cmd_en),
      .addr(br_addr),
      .wr_data(br_wr_data),
      .data_mask(br_data_mask),
      .rd_data(br_rd_data),
      .rd_data_valid(br_rd_data_valid),

      // inferred PSRAM ports
      .O_psram_ck(O_psram_ck),
      .O_psram_ck_n(O_psram_ck_n),
      .IO_psram_dq(IO_psram_dq),
      .IO_psram_rwds(IO_psram_rwds),
      .O_psram_cs_n(O_psram_cs_n),
      .O_psram_reset_n(O_psram_reset_n)
  );

  localparam RAM_DEPTH_BITWIDTH = 21;

  // ----------------------------------------------------------
  // -- RAMIO
  // ----------------------------------------------------------
  reg ramio_enable;
  reg [1:0] ramio_write_type;
  reg [2:0] ramio_read_type;
  reg [31:0] ramio_address;
  reg [31:0] ramio_data_in;
  wire [31:0] ramio_data_out;
  wire ramio_data_out_ready;
  wire ramio_busy;
  reg [5:0] ramio_leds;

  RAMIO #(
      .RAM_DEPTH_BITWIDTH(RAM_DEPTH_BITWIDTH),
      .RAM_ADDRESSING_MODE(0),  // addressing 8 bit words
      .CACHE_LINE_IX_BITWIDTH(5),
      .CLK_FREQ(20_250_000),
      .BAUD_RATE(9_600)
  ) ramio (
      .rst_n(sys_rst_n && rpll_lock && br_init_calib),
      .clk(br_clk_out),
      .enable(ramio_enable),
      .write_type(ramio_write_type),
      .read_type(ramio_read_type),
      .address(ramio_address),
      .data_in(ramio_data_in),
      .data_out(ramio_data_out),
      .data_out_ready(ramio_data_out_ready),
      .busy(ramio_busy),
      .leds(ramio_leds),
      .uart_tx(uart_tx),
      .uart_rx(uart_rx),

      // burst RAM wiring; prefix 'br_'
      .br_cmd(br_cmd),  // 0: read, 1: write
      .br_cmd_en(br_cmd_en),  // 1: cmd and addr is valid
      .br_addr(br_addr),  // see 'RAM_ADDRESSING_MODE'
      .br_wr_data(br_wr_data),  // data to write
      .br_data_mask(br_data_mask),  // always 0 meaning write all bytes
      .br_rd_data(br_rd_data),  // data out
      .br_rd_data_valid(br_rd_data_valid)  // rd_data is valid
  );

  // ----------------------------------------------------------
  localparam STARTUP_WAIT = 1_000_000;

  // localparam FLASH_TRANSFER_BYTES_NUM = 32'h0020_0000;
  localparam FLASH_TRANSFER_BYTES_NUM = 32'h0010_0000;

  // used while reading flash
  reg [23:0] flash_data_to_send;
  reg [4:0] flash_bits_to_send;
  reg [31:0] flash_counter;
  reg [7:0] flash_current_byte_out;
  reg [7:0] flash_current_byte_num;
  reg [7:0] flash_data_in[4];

  // used while reading flash to increment 'cache_address'
  reg [31:0] ramio_address_next;

  localparam STATE_INIT_POWER = 0;
  localparam STATE_LOAD_CMD_TO_SEND = 1;
  localparam STATE_SEND = 2;
  localparam STATE_LOAD_ADDRESS_TO_SEND = 3;
  localparam STATE_READ_DATA = 4;
  localparam STATE_START_WRITE = 5;
  localparam STATE_WRITE = 6;
  localparam STATE_TEST_1 = 7;
  localparam STATE_TEST_2 = 8;
  localparam STATE_DONE = 9;

  reg [4:0] state = 0;
  reg [4:0] return_state = 0;

  always_ff @(posedge br_clk_out, negedge sys_rst_n) begin
    if (!sys_rst_n || !rpll_lock || !br_init_calib) begin

      flash_counter <= 0;
      flash_clk <= 0;
      flash_mosi <= 0;
      flash_cs <= 1;

      ramio_enable <= 0;
      ramio_read_type <= 0;
      ramio_write_type <= 0;
      ramio_address <= 0;
      ramio_address_next <= 0;
      ramio_data_in <= 0;

      led[4:0] <= 5'b1_1111;

      state <= STATE_INIT_POWER;

    end else begin
      led[5] <= ~ramio_busy;

      case (state)

        STATE_INIT_POWER: begin
          if (flash_counter > STARTUP_WAIT) begin
            flash_counter <= 0;
            state <= STATE_LOAD_CMD_TO_SEND;
          end else begin
            flash_counter <= flash_counter + 1;
          end
        end

        STATE_LOAD_CMD_TO_SEND: begin
          flash_cs <= 0;
          flash_data_to_send[23-:8] <= 3;  // command 3: read
          flash_bits_to_send <= 8;
          state <= STATE_SEND;
          return_state <= STATE_LOAD_ADDRESS_TO_SEND;
        end

        STATE_LOAD_ADDRESS_TO_SEND: begin
          flash_data_to_send <= 0;  // address 0x0
          flash_bits_to_send <= 24;
          flash_current_byte_num <= 0;
          state <= STATE_SEND;
          return_state <= STATE_READ_DATA;
        end

        STATE_SEND: begin
          if (flash_counter == 0) begin
            // at clock to low
            flash_clk <= 0;
            flash_mosi <= flash_data_to_send[23];
            flash_data_to_send <= {flash_data_to_send[22:0], 1'b0};
            flash_bits_to_send <= flash_bits_to_send - 1;
            flash_counter <= 1;
          end else begin
            // at clock to high
            flash_counter <= 0;
            flash_clk <= 1;
            if (flash_bits_to_send == 0) begin
              state <= return_state;
            end
          end
        end

        STATE_READ_DATA: begin
          if (!flash_counter[0]) begin
            flash_clk <= 0;
            flash_counter <= flash_counter + 1;
            if (flash_counter[3:0] == 0 && flash_counter > 0) begin
              // every 16 clock ticks (8 bit * 2)
              flash_data_in[flash_current_byte_num] <= flash_current_byte_out;
              flash_current_byte_num <= flash_current_byte_num + 1;
              if (flash_current_byte_num == 3) begin
                state <= STATE_START_WRITE;
              end
            end
          end else begin
            flash_clk <= 1;
            flash_current_byte_out <= {flash_current_byte_out[6:0], flash_miso};
            flash_counter <= flash_counter + 1;
          end
        end

        STATE_START_WRITE: begin
          if (!ramio_busy) begin
            ramio_enable <= 1;
            ramio_read_type <= 0;
            ramio_write_type <= 2'b11;
            ramio_address <= ramio_address_next;
            ramio_address_next <= ramio_address_next + 4;
            ramio_data_in <= {
              flash_data_in[3], flash_data_in[2], flash_data_in[1], flash_data_in[0]
            };
            state <= STATE_WRITE;
          end
        end

        STATE_WRITE: begin
          if (!ramio_busy) begin
            ramio_enable <= 0;
            flash_current_byte_num <= 0;
            if (ramio_address_next < FLASH_TRANSFER_BYTES_NUM) begin
              state <= STATE_READ_DATA;
            end else begin
              flash_cs <= 1;
              state <= STATE_TEST_1;
            end
          end
        end

        STATE_TEST_1: begin
          if (!ramio_busy) begin
            // read unsigned half-word (16 bits) from address 0x4
            ramio_enable <= 1;
            ramio_read_type <= 3'b010;
            ramio_write_type <= 0;
            ramio_address <= 4;
            state <= STATE_TEST_2;
          end
        end

        STATE_TEST_2: begin
          if (ramio_data_out_ready) begin
            if (ramio_data_out == 32'h00_00_41_20) begin  // addr: 0x4, half-word
              led[4:0] <= 5'b0_0000;
            end else begin
              led[4:0] <= 5'b1_1110;
            end
            state <= STATE_DONE;
          end
        end

        STATE_DONE: begin
        end

      endcase
    end
  end

endmodule

`default_nettype wire
